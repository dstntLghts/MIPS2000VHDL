----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:45:14 09/26/2013 
-- Design Name: 
-- Module Name:    rom - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;


entity rom is 
port ( address  : in std_logic_vector (6 downto 0) ;
       data : out std_logic_vector( 63 downto 0 )
		 ) ;
end entity ;

------------------
architecture arch of rom is 
type memory is array ( 0 to 87 ) of std_logic_vector( 63 downto 0 ) ;
constant my_rom : memory := (
0  => "0100001000001110001001001000000000000000000001100000000000000100",
1  => "0100110110110101001001001001000010111001010111000000000000000111",
2  => "0111110101000100000001001110000010001111010100101000011000001000",
3  => "0010010110110000001001000001000011010001111011000000000010110010",
4  => "1000001000110101000001000001000010000000000000000000011000000000",
5  => "0101000001000110001001001111011010010001111000000000000000000100",
6  => "0100000001001000110101110111011011101000000000000000000000000000",
7  => "1100000000000001001001111111111000000000000000000000011011011000",
8  => "0110001100111000111001000011010011011010011010101001110111101000",
9  => "0101001000101001000001001000000000010000000000000000010000100100",
10 => "0101010000001110101001001001000010011010000000000000000011000000",
11 => "0100001000000010010011010110010100000001111100000100010000100100",
12 => "0000000101011011010001000101000001001000000000101100011111100001",
13 => "0111100001000110001000000001000001110010000000000000000110000010",
14 => "1010000111110101001001001000000011010001111000000000000000100000",
15 => "1010001101001100001110000001000000001101001101010000000000110010",
16 => "1100000001000001001000001111001100000000000000000000000001100100",
17 => "0000010010001010010010000000100000111001101001111100110110110001",
18 => "0000001000110101001001001001001011100000000000000000001100000000",
19 => "0101001001001001001001111111010100000110010010001000000001111001",
20 => "0001100110100001000001110001000010111011101000000011000000001000",
21 => "0001001000000000000001000001110111000000000000000000000000000001",
22 => "0000110001000001001000000010010100000000100000000011100000000000",
23 => "0001100111000111000101000101000011010011010101001110000010000101",
24 => "1111010100001000000001001000100000111101000110101100000000000100",
25 => "1001111000001001000101000000000000011100000000000001001011001000",
26 => "0100001000001110001001001001000100000000000000110000000000000100",
27 => "0101000000001001001110101001000000101010000000000110000000000000",
28 => "1110000001111100001011001011111110000000100011001011001111100110",
29 => "1010000110011100011100100001001000111101001101010100111010110010",
30 => "0001011101110001001001001110000001010110010000100000110000000010",
31 => "0100100101000101101100110100000100000011000000011100100111010110",
32 => "0100110101010111010100001001000000111110111110010011000010110010",
33 => "1011101001001000001001001000000010010000000000000000000000000011",
34 => "1000001000000001000110101000000011000000000011000000000000000000",
35 => "1111001001000001000001110010111100000000000011110001101111001001",
36 => "0100001001001000000000000110000100110000000000000000000000000100",
37 => "0010001100001000001000000110000010001010000011000000000000001000",
38 => "0111101001000000000000001000110011010011100000000000000000000100",
39 => "0101001001000000000101000001100100000000000001010100111110010010",
40 => "1111001001001001001001110011011000000000100000000111010000111111",
41 => "1000100101100101000101000001000010111111111010000000000010000101",
42 => "1000001111100001011000000000000001111111000100110100000000000100",
43 => "0100110001001000001001000110011000000000000000000001101001100000",
44 => "0000001000001001110100110111111000011000000000000000000000000100",
45 => "0101001000110000001001110110010100000000001101000000000001111111",
46 => "1110000010011101010010000011111110001010111100100111100001001001",
47 => "0000100111000010110000100111110001010101100011111101001010100101",
48 => "0100110001000001000110010010111000100000000011100000000001111111",
49 => "0010001111100001001001000101000000100100011001011000001000010010",
50 => "1001001110000001000001001000000001000000000000000000000001100100",
51 => "0001001000110100110010010011010100111000000000000000000101110100",
52 => "0010101010001111001000001000001000110010110100000000000000001100",
53 => "1001001000001001001000110101001011000000000110000000000000000000",
54 => "1100001000101001001001001001000011111011110000000000000000000111",
55 => "1011000100111010100001001000001010111101111001001100000010110010",
56 => "1001000111110000101100110001000010010010001100101100111000111010",
57 => "1110001111001110011010110110111001000001110100100000100100011001",
58 => "1001111101000100010110010011111100100111110110101111111011001111",
59 => "0100001001111011110110011111110101000000000000111000111000110010",
60 => "0001001011011000110100100001000001101000111101101001000000000001",
61 => "0100000000001001000110101000000010000000000110000000000000000000",
62 => "0100000001001000010111111111001100000100000000000000100100000111",
63 => "0101000001001110000010111111111101100100000000000000000001111101",
64 => "0100101001000001000000000110001010000000000000000000000010110100",
65 => "0101001000000001001001001000110001110000000000000000000000010000",
66 => "0000110011010001001000110001001001011101110110100000000110000010",
67 => "0101001001001001001001001001000100000000000000000000000000010101",
68 => "0001000000110001001001110010010110010001111000000000000000000100",
69 => "0001010001101001100000000000100011100001101001101000010000000000",
70 => "0100000110000001111110011111011100100001101100000000011100110111",
71 => "0111000001000001110001000000000010000010000000000000110000000010",
72 => "1000010100011010011100001000000010111000011010011010100000000100",
73 => "0000101100001000000001001001110000010001111110000000000000000010",
74 => "1111001000110001001001001001001000101100000000000000000000001001",
75 => "0000000111000000001000001111010000000000000001111000000000000100",
76 => "0011111101010001000000011110100111100011110101001010000000001110",
77 => "0100001000001110000001001001100000000000000110000000000000000000",
78 => "0100000110001111111000101101110010000000000000000011001101101000",
79 => "1001000000000001110101000000000010000000000000001100000000000000",
80 => "1100001011011000001110000000000001110011000011000000000011001000",
81 => "0110101000000001000000000001000100000000000000000001100000001000",
82 => "0100001001001001000001110001000100000001100000000000000000000001",
83 => "1001000001000110001000001001000001000000000000000011000000000001",
84 => "0000101001000000000000001000001010000000000000000000000000001000",
85 => "0011010010011000101000001110100011000010101100101000011000000000",
86 => "1001101001001100011101010110001011100001010110010100110001110001",
87 => "0100001000001000110000001000100000000000110000000000000000000100"
);
begin
   process (address)
   begin
     case address is
       when "0000000" => data <= my_rom(0);
       when "0000001" => data <= my_rom(1);
       when "0000010" => data <= my_rom(2);
       when "0000011" => data <= my_rom(3);
       when "0000100" => data <= my_rom(4);
       when "0000101" => data <= my_rom(5);
       when "0000110" => data <= my_rom(6);
       when "0000111" => data <= my_rom(7);
       when "0001000" => data <= my_rom(8);
       when "0001001" => data <= my_rom(9);
       when "0001010" => data <= my_rom(10);
       when "0001011" => data <= my_rom(11);
       when "0001100" => data <= my_rom(12);
       when "0001101" => data <= my_rom(13);
       when "0001110" => data <= my_rom(14);
       when "0001111" => data <= my_rom(15);		 
		 when "0010000" => data <= my_rom(16);
       when "0010001" => data <= my_rom(17);
       when "0010010" => data <= my_rom(18);
       when "0010011" => data <= my_rom(19);
       when "0010100" => data <= my_rom(20);
       when "0010101" => data <= my_rom(21);
       when "0010110" => data <= my_rom(22);
       when "0010111" => data <= my_rom(23);
       when "0011000" => data <= my_rom(24);
       when "0011001" => data <= my_rom(25);
       when "0011010" => data <= my_rom(26);
       when "0011011" => data <= my_rom(27);
       when "0011100" => data <= my_rom(28);
       when "0011101" => data <= my_rom(29);
       when "0011110" => data <= my_rom(30);
       when "0011111" => data <= my_rom(31);	 
		 when "0100000" => data <= my_rom(32);
       when "0100001" => data <= my_rom(33);
       when "0100010" => data <= my_rom(34);
       when "0100011" => data <= my_rom(35);
       when "0100100" => data <= my_rom(36);
       when "0100101" => data <= my_rom(37);
       when "0100110" => data <= my_rom(38);
       when "0100111" => data <= my_rom(39);
       when "0101000" => data <= my_rom(40);
       when "0101001" => data <= my_rom(41);
       when "0101010" => data <= my_rom(42);
       when "0101011" => data <= my_rom(43);
       when "0101100" => data <= my_rom(44);
       when "0101101" => data <= my_rom(45);
       when "0101110" => data <= my_rom(46);
       when "0101111" => data <= my_rom(47);		 
		 when "0110000" => data <= my_rom(48);
       when "0110001" => data <= my_rom(49);
       when "0110010" => data <= my_rom(50);
       when "0110011" => data <= my_rom(51);
       when "0110100" => data <= my_rom(52);
       when "0110101" => data <= my_rom(53);
       when "0110110" => data <= my_rom(54);
       when "0110111" => data <= my_rom(55);
       when "0111000" => data <= my_rom(56);
       when "0111001" => data <= my_rom(57);
       when "0111010" => data <= my_rom(58);
       when "0111011" => data <= my_rom(59);
       when "0111100" => data <= my_rom(60);
       when "0111101" => data <= my_rom(61);
       when "0111110" => data <= my_rom(62);
       when "0111111" => data <= my_rom(63);	 
		 when "1000000" => data <= my_rom(64);
       when "1000001" => data <= my_rom(65);
       when "1000010" => data <= my_rom(66);
       when "1000011" => data <= my_rom(67);
       when "1000100" => data <= my_rom(68);
       when "1000101" => data <= my_rom(69);
       when "1000110" => data <= my_rom(70);
       when "1000111" => data <= my_rom(71);
       when "1001000" => data <= my_rom(72);
       when "1001001" => data <= my_rom(73);
       when "1001010" => data <= my_rom(74);
       when "1001011" => data <= my_rom(75);
       when "1001100" => data <= my_rom(76);
       when "1001101" => data <= my_rom(77);
       when "1001110" => data <= my_rom(78);
       when "1001111" => data <= my_rom(79);		 
		 when "1010000" => data <= my_rom(80);
       when "1010001" => data <= my_rom(81);
       when "1010010" => data <= my_rom(82);
       when "1010011" => data <= my_rom(83);
       when "1010100" => data <= my_rom(84);
       when "1010101" => data <= my_rom(85);
       when "1010110" => data <= my_rom(86);
       when "1010111" => data <= my_rom(87);
       when others => data <= x"0000000000000000";
	 end case;
  end process;
end arch;